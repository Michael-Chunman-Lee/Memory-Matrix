module MemoryMatrix(
	input CLOCK_50);
endmodule